//module LAB2(a,b,c,d,e,f,g,h,i,j,k);   
//      input a,b,c,d;
//      output e,f,g,h,i,j,k;
//      assign e = ((~a & ~b & ~c & d) | (~a & b & ~c & ~d) | (a & ~b & c & d) | (a & b & ~c & d));
//      assign f = ((~a & b & ~c & d) | (~a & b & c & ~d) | (a & ~b & c & d) | (a & b & ~c & ~d) | (a & b & c & ~d) | (a & b & c & d));
//      assign g = ((~a & ~b & c & ~d) | (a & b & ~c & ~d) | (a & b & c & ~d) | (a & b & c & d));
//      assign h = ((~a & ~b & ~c & d) | (~a & b & ~c & ~d) | (~a & b & c & d) | (a & ~b & c & ~d) | (a & b & c & d));
//      assign i = ((~a & ~b & ~c & d) | (~a & ~b & c & d) | (~a & b & ~c & ~d) | (~a & b & ~c & d) | (~a & b & c & d) | (a & ~b & ~c & d));
//      assign j = ((~a & ~b & ~c & d) | (~a & ~b & c & ~d) | (~a & ~b & c & d) | (~a & b & c & d) | (a & b & ~c & d));
//      assign k = ((~a & ~b & ~c & ~d) | (~a & ~b & ~c & d) | (~a & b & c & d) | (a & b & ~c & ~d)); 
//endmodule

module LAB2(a,b);
input [3:0] a;
output [6:0] b;

assign b[0] = ((~a[3] & ~a[2] & ~a[1] & a[0]) | (~a[3] & a[2] & ~a[1] & ~a[0]) | (a[3] & ~a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & a[0]));
assign b[1] = ((~a[3] & a[2] & ~a[1] & a[0]) | (~a[3] & a[2] & a[1] & ~a[0]) | (a[3] & ~a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & ~a[0]) | (a[3] & a[2] & a[1] & ~a[0]) | (a[3] & a[2] & a[1] & a[0]));
assign b[2] = ((~a[3] & ~a[2] & a[1] & ~a[0]) | (a[3] & a[2] & ~a[1] & ~a[0]) | (a[3] & a[2] & a[1] & ~a[0]) | (a[3] & a[2] & a[1] & a[0]));
//assign b[2] = ((~a[3] & ~a[2] & a[1] & ~a[0]) | (a[3] & a[1] & ~a[0]) | (a[2] & a[1] & a[0]));
assign b[3] = ((~a[3] & ~a[2] & ~a[1] & a[0]) | (~a[3] & a[2] & ~a[1] & ~a[0]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & ~a[2] & a[1] & ~a[0]) | (a[3] & a[2] & a[1] & a[0]));
assign b[4] = ((~a[3] & ~a[2] & ~a[1] & a[0]) | (~a[3] & ~a[2] & a[1] & a[0]) | (~a[3] & a[2] & ~a[1] & ~a[0]) | (~a[3] & a[2] & ~a[1] & a[0]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & ~a[2] & ~a[1] & a[0]));
assign b[5] = ((~a[3] & ~a[2] & ~a[1] & a[0]) | (~a[3] & ~a[2] & a[1] & ~a[0]) | (~a[3] & ~a[2] & a[1] & a[0]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & a[0]));
//assign b[6] = ((~a[3] & ~a[2] & ~a[1] & ~a[0]) | (~a[3] & ~a[2] & ~a[1] & a[0]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & ~a[0]));
assign b[6] = ((~a[3] & ~a[2] & ~a[1]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & ~a[0]));
 
endmodule

//part 3

//assign b[6] = ((~a[3] & ~a[2] & ~a[1]) | (~a[3] & a[2] & a[1] & a[0]) | (a[3] & a[2] & ~a[1] & ~a[0]));